// Binary to gray converter

module Binary_to_Gray_Converter #(
  parameter VEC_W = 4
)(
  input     wire[VEC_W-1:0] bin_i,
  output    wire[VEC_W-1:0] gray_o // update all functions !!

);

  
endmodule